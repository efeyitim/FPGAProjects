-------------------------------------------------------------------------------
-- Title      : Testbench for design "multiplicator"
-- Project    : 
-------------------------------------------------------------------------------
-- File	      : multiplicator_tb.vhd
-- Author     : Efe  <efe@efeASUS>
-- Company    : 
-- Created    : 2022-07-15
-- Last update: 2022-07-15
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2022 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date	       Version	Author	Description
-- 2022-07-15  1.0	efe	Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------

entity multiplicator_tb is

end entity multiplicator_tb;

--------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------

architecture tb of multiplicator_tb is

    -- component generics
    constant LENGTH : integer := 5;

    -- component ports
    signal clk		: std_logic := '0';
    signal rst_n	: std_logic;
    signal en		: std_logic;
    signal multiplicand : std_logic_vector(2**LENGTH-1 downto 0);
    signal multiplier	: std_logic_vector(2**LENGTH-1 downto 0);
    signal product	: std_logic_vector(2**(LENGTH+1)-1 downto 0);
    signal busy		: std_logic;
    signal done		: std_logic;


begin  -- architecture tb

    -- component instantiation
    DUT : entity work.multiplicator
	generic map (
	    LENGTH	 => LENGTH)
	port map (
	    clk		 => clk,
	    rst_n	 => rst_n,
	    en		 => en,
	    multiplicand => multiplicand,
	    multiplier	 => multiplier,
	    product	 => product,
	    busy	 => busy,
	    done	 => done);

    -- clock generation
    clk <= not clk after 10 ns;

    PROC_TB		: process is
	constant period : time := 20 ns;
    begin  -- process PROC_TB
	rst_n		       <= '0';
	en		       <= '0';
	multiplicand	       <= (others => '0');
	multiplier	       <= (others => '0');
	wait for 5*period;
	rst_n		       <= '1';
	wait for 5*period;
	multiplicand	       <= x"00000017";
	multiplier	       <= x"00000013";
	wait for 5*period;
	en		       <= '1';
	wait for period;
	en		       <= '0';
	wait for period;
	en		       <= '1';
	multiplicand	       <= x"0000000B";
	multiplier	       <= x"00000003";
	wait for 35*period;
	en		       <= '0';
	wait on busy;
	multiplicand	       <= x"00010D48";	-- 68936d
	multiplier	       <= x"00001119";	-- 4377d, product = 301732872d = 11FC1408
	en		       <= '1';
	wait on busy;
	en		       <= '0';
	wait on busy;
	multiplicand	       <= x"FFFFCDB8";	-- -3248d
	multiplier	       <= x"0000F4DA";	-- 62682, product = 301732872d = ECABFC770
	en		       <= '1';
	wait on busy;
	en <= '0';
	wait on busy;
	multiplicand	       <= x"FFFFDF82";	-- -8318
	multiplier	       <= x"FFFFCEBA";	-- -12614, product = 06410074h
	en		       <= '1';
	wait on busy;
	en <= '0';
	wait on busy;	

	wait for 10 us;
    end process PROC_TB;
end architecture tb;
